module vxai

import json
import net.http

// The API path for completions.
pub const completion_path = 'completions'

// CompletionInput represents the input parameters for a completion request.
// It includes options for customizing the behavior and output of the model.
pub struct CompletionInput {
pub:
	// The prompt to generate completions for.
	prompt string

	// Number between -2.0 and 2.0. Positive values penalize new tokens based on
	// their existing frequency in the text so far, decreasing the model's
	// likelihood to repeat the same line verbatim.
	frequency_penalty ?f32

	// A JSON object that maps tokens (specified by their token ID in the tokenizer)
	// to an associated bias value from -100 to 100. Mathematically, the bias is added
	// to the logits generated by the model prior to sampling. The exact effect will
	// vary per model, but values between -1 and 1 should decrease or increase likelihood
	// of selection; values like -100 or 100 should result in a ban or exclusive selection
	//  of the relevant token.
	logit_bias ?map[string]f32

	// Whether to return log probabilities of the output tokens or not. If true, returns
	// the log probabilities of each output token returned in the content of message.
	logprobs ?bool

	// The maximum number of tokens that can be generated in the chat completion. This
	// value can be used to control costs for text generated via API.
	max_tokens ?int

	// Specifies the model to be used for the request.
	model string

	// How many chat completion choices to generate for each input message. Note that
	// you will be charged based on the number of generated tokens across all of the
	// choices. Keep n as 1 to minimize costs.
	n ?int

	// Number between -2.0 and 2.0. Positive values penalize new tokens based on whether
	// they appear in the text so far, increasing the model's likelihood to talk about new topics.
	presence_penalty ?f32

	// response_format specifies the format of the response, such as plain text or JSON.
	// When null, the default format is used.
	response_format ?string

	// If specified, our system will make a best effort to sample deterministically, such that
	// repeated requests with the same `seed` and parameters should return the same result.
	// Determinism is not guaranteed, and you should refer to the `system_fingerprint` response
	// parameter to monitor changes in the backend.
	seed ?int

	// Up to 4 sequences where the API will stop generating further tokens.
	stop ?[]string

pub mut:
	// If set, partial message deltas will be sent. Tokens will be sent as data-only server-sent
	// events as they become available, with the stream terminated by a `data: [DONE]` message.
	stream bool

	// What sampling temperature to use, between 0 and 2. Higher values like 0.8 will make the
	// output more random, while lower values like 0.2 will make it more focused and deterministic.
	temperature ?f32

	// An alternative to sampling with temperature, called nucleus sampling, where the model
	// considers the results of the tokens with top_p probability mass. So 0.1 means only the
	// tokens comprising the top 10% probability mass are considered. It is generally recommended
	// to alter this or `temperature` but not both.
	top_p ?f32

	// A unique identifier representing your end-user, which can help xAI to monitor and detect abuse
	user ?string

}

// CompletionInput.new creates a new CompletionInput instance with the given prompt and model.
//
// Parameters:
// - prompt: The input text to generate a completion for.
// - model: The name of the model to use for generating the completion.
//
// Returns:
// - A new CompletionInput instance.
pub fn CompletionInput.new(prompt string, model string) CompletionInput {
	return CompletionInput{
		prompt: prompt
		model:  model
	}
}

// CompletionResponse represents the response from a text completion API call.
// It includes the generated choices, metadata about the request, and token usage details.
pub struct CompletionResponse {
pub:
	// choices contains the list of generated completions.
	choices []CompletionChoice

	// created is the Unix timestamp indicating when the response was generated.
	created i64

	// id is a unique identifier for this completion response.
	id string

	// model specifies the model used to generate the completion.
	model string

	// object specifies the type of object returned, typically "text_completion".
	object string

	// system_fingerprint is a server-generated identifier for debugging or tracking.
	system_fingerprint string

	// usage provides token usage details, including prompt and completion token counts.
	usage CompletionUsage
}

// CompletionChoice represents an individual generated completion within the response.
pub struct CompletionChoice {
pub:
	// finish_reason indicates why the generation stopped (e.g., "length", "stop").
	finish_reason string

	// index is the position of this choice in the list of returned choices.
	index int

	// text contains the generated text for this completion.
	text string
}

// CompletionUsage provides statistics on token usage for a completion request.
pub struct CompletionUsage {
pub:
	// completion_tokens is the number of tokens in the generated completion.
	completion_tokens int

	// prompt_tokens is the number of tokens in the input prompt.
	prompt_tokens int

	// total_tokens is the total number of tokens processed (prompt + completion).
	total_tokens int
}

// StreamCompletionChunk represents a single streamed chunk of a completion response.
pub struct StreamCompletionChunk {
pub:
	// id is a unique identifier for this specific chunk of the completion.
	id string

	// object specifies the type of the returned object, typically "completion.chunk".
	object string

	// created is the Unix timestamp (in seconds) indicating when this chunk was generated.
	created i64

	// choices is an array of StreamCompletionChoice objects, each representing a portion of the streamed completion.
	choices []StreamCompletionChoice

	// usage contains token usage statistics for this chunk, including prompt and completion tokens.
	usage StreamCompletionUsage

	// system_fingerprint is a server-generated identifier for debugging or reference.
	system_fingerprint string
}

// StreamCompletionChoice represents an individual choice within a streamed chunk.
pub struct StreamCompletionChoice {
pub:
	// index is the position of this choice in the list of returned choices.
	index int

	// delta contains newly streamed content or role information for this choice.
	delta StreamCompletionDelta

	// finish_reason is an optional reason indicating why this choice concluded (e.g., "stop").
	finish_reason ?string
}

// StreamCompletionUsage contains token usage details for a streamed completion segment.
pub struct StreamCompletionUsage {
pub:
	// prompt_tokens is the number of tokens used in the input prompt.
	prompt_tokens int

	// completion_tokens is the number of tokens generated in this streamed response.
	completion_tokens int

	// total_tokens is the total number of tokens processed so far (prompt + completion).
	total_tokens int

	// prompt_tokens_details provides a detailed breakdown of the input tokens by type (e.g., text, audio).
	prompt_tokens_details StreamCompletionPromptTokenDetails
}

// StreamCompletionPromptTokenDetails provides a breakdown of the prompt tokens by type.
pub struct StreamCompletionPromptTokenDetails {
pub:
	// text_tokens is the number of tokens derived from textual input.
	text_tokens int

	// audio_tokens is the number of tokens derived from audio input.
	audio_tokens int

	// image_tokens is the number of tokens derived from image input.
	image_tokens int

	// cached_tokens is the number of tokens retrieved from cache.
	cached_tokens int
}

// StreamCompletionDelta represents incremental updates to the streamed completion.
pub struct StreamCompletionDelta {
pub:
	// content is the newly generated text or partial completion content, if any.
	content ?string

	// role is the role associated with this content, such as "assistant" or "system".
	role string
}

// get_completion sends a completion request to the API.
//
// Parameters:
// - input: A CompletionInput instance containing the request parameters.
//
// Returns:
// - A CompletionResponse containing the generated completions.
// - An error if the request fails or if the response cannot be decoded.
pub fn (c XAIClient) get_completion(input CompletionInput) !CompletionResponse {
	data := json.encode(input)
	res := c.post(vxai.completion_path, data) or { return error('Failed to post completion') }
	return json.decode(CompletionResponse, res.body) or { return err }
}

// stream_completion sends a streaming completion request to the API.
//
// Parameters:
// - input: A mutable CompletionInput instance containing the request parameters.
// - on_message: A callback function invoked for each streamed chunk of the completion.
// - on_finish: A callback function invoked when streaming finishes.
//
// Returns:
// - An HTTP response object for the streaming request.
// - An error if the request fails.
pub fn (c XAIClient) stream_completion(mut input CompletionInput, on_message fn (StreamOnMessageFn), on_finish fn ()) !http.Response {
	input.stream = true
	data := json.encode(input)
	return c.stream(vxai.completion_path, data, on_message, on_finish) or { return err }
}
