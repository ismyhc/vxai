module vxai

import json
import net.http

// ChatCompletionInput represents the input structure for creating a chat completion.
// It contains various parameters to control the behavior and output of the model.
pub struct ChatCompletionInput {
pub:
	// frequency_penalty adjusts the likelihood of repetitive token generation.
	// A higher value discourages repetition in the response.
	frequency_penalty ?f32

	// logit_bias allows specific tokens to be biased by modifying their logits.
	// It maps tokens (strings) to their respective bias values.
	logit_bias ?map[string]f32

	// logprobs specifies whether to include the log probabilities of tokens in the response.
	// When true, the response will contain token-level probabilities.
	logprobs ?bool

	// max_tokens sets the maximum number of tokens the model can generate.
	// This limits the length of the output.
	max_tokens ?int

	// messages contains the conversation history as an array of ChatCompletionMessage.
	// It provides context for the assistant to generate appropriate responses.
	messages []ChatCompletionMessage

	// model specifies the name of the model to use for the chat completion.
	// This determines the capabilities and behavior of the assistant.
	model string

	// n defines the number of completions to generate.
	// For example, setting n=2 will produce two independent responses.
	n ?int

	// presence_penalty adjusts the likelihood of introducing new topics in the response.
	// A higher value encourages diverse and novel content.
	presence_penalty ?f32

	// response_format specifies the format of the response, such as plain text or JSON.
	// When null, the default format is used.
	response_format ?string

	// seed sets the random seed for reproducibility.
	// Using the same seed produces consistent results for the same input.
	seed ?int

	// stop defines sequences where the model should stop generating text.
	// This prevents the model from continuing beyond certain keywords or phrases.
	stop ?[]string

	// stream enables or disables response streaming.
	// When true, the response is sent as a stream rather than a complete object.
	stream bool

	// temperature controls the randomness of the response generation.
	// A lower value makes the output more focused, while a higher value makes it more creative.
	temperature ?f32

	// tool_choice specifies the tool the model should use for generating the response.
	// This allows fine-grained control over the assistant's behavior.
	tool_choice ?string

	// tools lists the tools available for the model to use.
	// For example, it could include summarization or translation tools.
	tools ?[]string

	// top_logprobs sets the number of top tokens to return log probabilities for.
	// This is useful for inspecting token-level probabilities.
	top_logprobs ?int

	// top_p enables nucleus sampling, limiting the probability space to the top p percentage.
	// This controls the diversity of the response.
	top_p ?f32

	// user identifies the end user of the request.
	// This can be used for analytics or personalization.
	user ?string
}

// ChatCompletionMessage represents a message exchanged during a chat completion.
// Each message has a role and its corresponding content.
pub struct ChatCompletionMessage {
pub:
	// role specifies the role of the message sender.
	// Examples include "user", "assistant", or "system".
	role string

	// content contains the text of the message.
	// This is the actual message exchanged in the conversation.
	content string
}

// Choice represents an individual choice or completion generated by the model.
// It includes information about the generated message and its metadata.
pub struct Choice {
pub:
	// finish_reason indicates why the completion ended.
	// Examples include "stop" (end of generation) or "length" (max tokens reached).
	finish_reason string

	// index is the position of this choice in the list of completions.
	index int

	// message is the generated message for this choice.
	// It contains the content and role of the response.
	message ChatCompletionMessage
}

// Usage provides details about token usage for a chat completion request.
// It includes counts for prompt, completion, and total tokens.
pub struct Usage {
pub:
	// completion_tokens is the number of tokens used in the generated response.
	completion_tokens int

	// prompt_tokens is the number of tokens used in the input prompt.
	prompt_tokens int

	// total_tokens is the total number of tokens used in the request and response.
	// This is the sum of completion_tokens and prompt_tokens.
	total_tokens int
}

// ChatCompletionResponse represents the response from the chat completion API.
// It includes the generated choices, metadata, and token usage information.
pub struct ChatCompletionResponse {
pub:
	// choices is a list of choices generated by the model.
	// Each choice includes a generated message and its associated metadata.
	choices []Choice

	// created is a Unix timestamp indicating when the response was created.
	created i64

	// id is a unique identifier for the response.
	id string

	// model specifies the name of the model used for the chat completion.
	model string

	// object is the type of object represented by this response.
	// Typically, this is "chat.completion".
	object string

	// system_fingerprint is a unique fingerprint for the system handling the request.
	system_fingerprint string

	// usage provides details about the token usage for the request and response.
	usage Usage
}

// StreamChatCompletionChunk represents a single streamed chunk of a chat completion response.
pub struct StreamChatCompletionChunk {
pub:
	// A unique identifier for this specific chunk of the completion.
	id string
	// The type of the returned object, typically "chat.completion.chunk".
	object string
	// The Unix timestamp (in seconds) indicating when this chunk was generated.
	created i64
	// An array of StreamChoice objects, each representing a portion of the streamed completion.
	choices []StreamChoice
	// Token usage statistics for this chunk, including prompt and completion tokens.
	usage StreamUsage
	// A server-generated fingerprint for debugging or reference.
	system_fingerprint string
}

// StreamChoice represents an individual choice within a streamed chunk.
pub struct StreamChoice {
pub:
	// The position of this choice in the list of returned choices.
	index int
	// A StreamDelta object containing newly streamed content or role information.
	delta StreamDelta
	// An optional reason indicating why this choice concluded (e.g., "stop").
	finish_reason ?string
}

// StreamUsage contains token usage details for a streamed completion segment.
pub struct StreamUsage {
pub:
	// The number of tokens used in the prompt.
	prompt_tokens int
	// The number of tokens generated in this streamed response.
	completion_tokens int
	// The total number of tokens processed so far (prompt + completion).
	total_tokens int
	// Detailed breakdown of the prompt tokens by type (text, audio, image, cached).
	prompt_tokens_details PromptTokenDetails
}

// PromptTokenDetails provides a breakdown of the prompt tokens by type.
pub struct PromptTokenDetails {
pub:
	// Number of tokens derived from textual input.
	text_tokens int
	// Number of tokens derived from audio input.
	audio_tokens int
	// Number of tokens derived from images.
	image_tokens int
	// Number of tokens retrieved from cache.
	cached_tokens int
}

// StreamDelta represents incremental updates to the streamed completion.
pub struct StreamDelta {
pub:
	// Newly generated text or partial completion content (if any).
	content ?string
	// The role associated with this content, such as "assistant" or "system".
	role string
}

// new creates a new instance of ChatCompletionInput.
//
// Parameters:
// - messages: A list of ChatCompletionMessage objects representing the conversation history.
// - model: The name of the model to use for generating the chat completion.
//
// Returns:
// - A new instance of ChatCompletionInput.
pub fn ChatCompletionInput.new(messages []ChatCompletionMessage, model string) ChatCompletionInput {
	return ChatCompletionInput{
		messages: messages
		model:    model
		stream:   true
	}
}

// get_chat_completion sends a chat completion request to the X.AI API and retrieves the response.
//
// Parameters:
// - input: A ChatCompletionInput struct containing the messages and model information for the request.
//
// Returns:
// - A ChatCompletionResponse struct containing the generated chat completion and metadata.
// - An error if the request fails or the response cannot be decoded.
pub fn (c XAIClient) get_chat_completion(input ChatCompletionInput) !ChatCompletionResponse {
	data := json.encode(input)
	res := c.post('chat/completions', data) or { return error('Failed to post chat completion') }
	return json.decode(ChatCompletionResponse, res.body) or { return err }
}

// stream_chat_completion sends a streaming chat completion request to the XAI API using the specified `input`.
//
// Each chunk of the streamed response is decoded as a `StreamChatCompletionChunk` and passed to the `on_message` callback
// as soon as it arrives. This allows you to process the streaming content incrementally rather than waiting for the full response.
//
// Parameters:
// - `input`: A `ChatCompletionInput` struct containing the details of the chat prompt and configuration for the completion.
// - `on_message`: A callback function of type `fn (StreamChatCompletionChunk)` that is invoked for each chunk of streamed data as it arrives.
//
// Returns:
// - `http.Response` representing the final HTTP response after the stream completes.
//
// Errors:
// Returns an error if the request fails to send, encounters connectivity issues, or if the response is invalid.
pub fn (c XAIClient) stream_chat_completion(input ChatCompletionInput, on_message fn (StreamChatCompletionChunk), on_finish fn ()) !http.Response {
	data := json.encode(input)
	return c.stream('chat/completions', data, on_message, on_finish) or { return err }
}
