module vxai

import json
import net.http

// The API path for chat completions.
pub const chat_completion_path = 'chat/completions'

// ChatCompletionInput represents the input parameters for a chat completion request.
// It includes options for customizing the behavior and output of the model.
pub struct ChatCompletionInput {
pub:
	// Number between -2.0 and 2.0. Positive values penalize new tokens based on
	// their existing frequency in the text so far, decreasing the model's
	// likelihood to repeat the same line verbatim.
	frequency_penalty ?f32

	// A JSON object that maps tokens (specified by their token ID in the tokenizer)
	// to an associated bias value from -100 to 100. Mathematically, the bias is added
	// to the logits generated by the model prior to sampling. The exact effect will
	// vary per model, but values between -1 and 1 should decrease or increase likelihood
	// of selection; values like -100 or 100 should result in a ban or exclusive selection
	//  of the relevant token.
	logit_bias ?map[string]f32

	// Whether to return log probabilities of the output tokens or not. If true, returns
	// the log probabilities of each output token returned in the content of message.
	logprobs ?bool

	// The maximum number of tokens that can be generated in the chat completion. This
	// value can be used to control costs for text generated via API.
	max_tokens ?int

	// A list of messages that make up the the chat conversation. Different models
	// support different message types, such as image and text.
	messages []ChatCompletionMessage

	// Model name for the model to use.
	model string

	// How many chat completion choices to generate for each input message. Note that
	// you will be charged based on the number of generated tokens across all of the
	// choices. Keep n as 1 to minimize costs.
	n ?int

	// Number between -2.0 and 2.0. Positive values penalize new tokens based on whether
	// they appear in the text so far, increasing the model's likelihood to talk about new topics.
	presence_penalty ?f32

	// response_format specifies the format of the response, such as plain text or JSON.
	// When null, the default format is used.
	response_format ?string

	// If specified, our system will make a best effort to sample deterministically, such that
	// repeated requests with the same `seed` and parameters should return the same result.
	// Determinism is not guaranteed, and you should refer to the `system_fingerprint` response
	// parameter to monitor changes in the backend.
	seed ?int

	// Up to 4 sequences where the API will stop generating further tokens.
	stop ?[]string

pub mut:
	// If set, partial message deltas will be sent. Tokens will be sent as data-only server-sent
	// events as they become available, with the stream terminated by a `data: [DONE]` message.
	stream bool

	// What sampling temperature to use, between 0 and 2. Higher values like 0.8 will make the
	// output more random, while lower values like 0.2 will make it more focused and deterministic.
	temperature ?f32

	// A list of tools the model may call. Currently, only functions are supported as a tool. Use
	// this to provide a list of functions the model may generate JSON inputs for. A max of 128
	// functions are supported.
	tool_choice ?string
	tools       ?[]string

	// An integer between 0 and 20 specifying the number of most likely tokens to return at each
	// token position, each with an associated log probability. logprobs must be set to true if
	// this parameter is used.
	top_logprobs ?int

	// An alternative to sampling with temperature, called nucleus sampling, where the model
	// considers the results of the tokens with top_p probability mass. So 0.1 means only the
	// tokens comprising the top 10% probability mass are considered. It is generally recommended
	// to alter this or `temperature` but not both.
	top_p ?f32

	// A unique identifier representing your end-user, which can help xAI to monitor and detect abuse
	user ?string

}

// ChatCompletionInput.new creates a new ChatCompletionInput with the given messages and model.
//
// Parameters:
// - messages: A list of input messages defining the conversation context.
// - model: The name of the model to use for the completion.
//
// Returns:
// - A ChatCompletionInput instance with the specified parameters.
pub fn ChatCompletionInput.new(messages []ChatCompletionMessage, model string) ChatCompletionInput {
	return ChatCompletionInput{
		messages: messages
		model:    model
	}
}

// ChatCompletionMessage represents a single message in the chat conversation.
pub struct ChatCompletionMessage {
pub:
	// role is the role of the message sender (e.g., "user", "assistant", "system").
	role string

	// content is the text content of the message.
	content string
}

// ChatCompletionChoice represents a single completion choice returned by the API.
pub struct ChatCompletionChoice {
pub:
	// finish_reason explains why the completion stopped (e.g., "length", "stop").
	finish_reason string

	// index is the position of this choice in the list of returned choices.
	index int

	// message contains the content of the generated message.
	message ChatCompletionMessage
}

// ChatCompletionUsage provides details about token usage for a request and response.
pub struct ChatCompletionUsage {
pub:
	// completion_tokens is the number of tokens in the generated response.
	completion_tokens int

	// prompt_tokens is the number of tokens in the input prompt.
	prompt_tokens int

	// total_tokens is the total number of tokens used (prompt + completion).
	total_tokens int
}

// ChatCompletionResponse represents the full response from the chat completion API.
pub struct ChatCompletionResponse {
pub:
	// choices contains the list of generated messages.
	choices []ChatCompletionChoice

	// created is the Unix timestamp when the response was generated.
	created i64

	// id is the unique identifier for this API response.
	id string

	// model specifies the model used for this completion.
	model string

	// object specifies the type of object returned (e.g., "text_completion").
	object string

	// system_fingerprint provides a system-level tracking identifier.
	system_fingerprint string

	// usage provides details about token usage in the request and response.
	usage ChatCompletionUsage
}

// StreamChatCompletionChunk represents a single chunk of a streamed response.
pub struct StreamChatCompletionChunk {
pub:
	// id is the unique identifier for this chunk.
	id string

	// object specifies the type of object returned.
	object string

	// created is the Unix timestamp when this chunk was generated.
	created i64

	// choices contains the partial completion choices in this chunk.
	choices []StreamChatCompletionChoice

	// usage provides token usage information for this chunk.
	usage StreamChatCompletionUsage

	// system_fingerprint provides a system-level tracking identifier for this chunk.
	system_fingerprint string
}

// StreamChatCompletionChoice represents a single partial completion returned during streaming.
pub struct StreamChatCompletionChoice {
pub:
	// index is the position of this choice in the list of streamed choices.
	index int

	// delta contains the incremental message content for this choice.
	delta StreamChatCompletionDelta

	// finish_reason explains why this choice's generation stopped (if applicable).
	finish_reason ?string
}

// StreamChatCompletionUsage provides token usage details for a streaming request.
pub struct StreamChatCompletionUsage {
pub:
	// prompt_tokens is the number of tokens in the input prompt.
	prompt_tokens int

	// completion_tokens is the number of tokens generated so far.
	completion_tokens int

	// total_tokens is the total number of tokens used (prompt + completion).
	total_tokens int

	// prompt_tokens_details provides a detailed breakdown of the input tokens.
	prompt_tokens_details StreamChatCompletionPromptTokenDetails
}

// StreamChatCompletionPromptTokenDetails provides a breakdown of tokens in the input prompt.
pub struct StreamChatCompletionPromptTokenDetails {
pub:
	// text_tokens is the number of tokens from text inputs.
	text_tokens int

	// audio_tokens is the number of tokens from audio inputs.
	audio_tokens int

	// image_tokens is the number of tokens from image inputs.
	image_tokens int

	// cached_tokens is the number of tokens retrieved from cache.
	cached_tokens int
}

// StreamChatCompletionDelta represents an incremental update to a message during streaming.
pub struct StreamChatCompletionDelta {
pub:
	// content is the partial message content for this update.
	content ?string

	// role is the role of the message sender for this update.
	role string
}

// get_chat_completion sends a chat completion request to the API.
//
// Parameters:
// - input: A ChatCompletionInput instance containing the request parameters.
//
// Returns:
// - A ChatCompletionResponse containing the generated completions.
// - An error if the request fails or if the response cannot be decoded.
pub fn (c XAIClient) get_chat_completion(input ChatCompletionInput) !ChatCompletionResponse {
	data := json.encode(input)
	res := c.post(vxai.chat_completion_path, data) or {
		return error('Failed to post chat completion')
	}
	return json.decode(ChatCompletionResponse, res.body) or { return err }
}

// stream_chat_completion sends a streaming chat completion request to the API.
//
// Parameters:
// - input: A mutable ChatCompletionInput instance containing the request parameters.
// - on_message: A callback function invoked for each streamed chunk.
// - on_finish: A callback function invoked when streaming finishes.
//
// Returns:
// - The HTTP response object for the streaming request.
// - An error if the request fails.
pub fn (c XAIClient) stream_chat_completion(mut input ChatCompletionInput, on_message fn (StreamOnMessageFn), on_finish fn ()) !http.Response {
	input.stream = true
	data := json.encode(input)
	return c.stream(vxai.chat_completion_path, data, on_message, on_finish) or { return err }
}
