module vxai

import json

// ChatCompletionInput represents the input structure for creating a chat completion.
// It contains various parameters to control the behavior and output of the model.
pub struct ChatCompletionInput {
pub:
	// frequency_penalty adjusts the likelihood of repetitive token generation.
	// A higher value discourages repetition in the response.
	frequency_penalty ?f32

	// logit_bias allows specific tokens to be biased by modifying their logits.
	// It maps tokens (strings) to their respective bias values.
	logit_bias ?map[string]f32

	// logprobs specifies whether to include the log probabilities of tokens in the response.
	// When true, the response will contain token-level probabilities.
	logprobs ?bool

	// max_tokens sets the maximum number of tokens the model can generate.
	// This limits the length of the output.
	max_tokens ?int

	// messages contains the conversation history as an array of ChatCompletionMessage.
	// It provides context for the assistant to generate appropriate responses.
	messages []ChatCompletionMessage

	// model specifies the name of the model to use for the chat completion.
	// This determines the capabilities and behavior of the assistant.
	model string

	// n defines the number of completions to generate.
	// For example, setting n=2 will produce two independent responses.
	n ?int

	// presence_penalty adjusts the likelihood of introducing new topics in the response.
	// A higher value encourages diverse and novel content.
	presence_penalty ?f32

	// response_format specifies the format of the response, such as plain text or JSON.
	// When null, the default format is used.
	response_format ?string

	// seed sets the random seed for reproducibility.
	// Using the same seed produces consistent results for the same input.
	seed ?int

	// stop defines sequences where the model should stop generating text.
	// This prevents the model from continuing beyond certain keywords or phrases.
	stop ?[]string

	// stream enables or disables response streaming.
	// When true, the response is sent as a stream rather than a complete object.
	stream bool

	// temperature controls the randomness of the response generation.
	// A lower value makes the output more focused, while a higher value makes it more creative.
	temperature ?f32

	// tool_choice specifies the tool the model should use for generating the response.
	// This allows fine-grained control over the assistant's behavior.
	tool_choice ?string

	// tools lists the tools available for the model to use.
	// For example, it could include summarization or translation tools.
	tools ?[]string

	// top_logprobs sets the number of top tokens to return log probabilities for.
	// This is useful for inspecting token-level probabilities.
	top_logprobs ?int

	// top_p enables nucleus sampling, limiting the probability space to the top p percentage.
	// This controls the diversity of the response.
	top_p ?f32

	// user identifies the end user of the request.
	// This can be used for analytics or personalization.
	user ?string
}

// ChatCompletionMessage represents a message exchanged during a chat completion.
// Each message has a role and its corresponding content.
pub struct ChatCompletionMessage {
pub:
	// role specifies the role of the message sender.
	// Examples include "user", "assistant", or "system".
	role string

	// content contains the text of the message.
	// This is the actual message exchanged in the conversation.
	content string
}

// Choice represents an individual choice or completion generated by the model.
// It includes information about the generated message and its metadata.
pub struct Choice {
pub:
	// finish_reason indicates why the completion ended.
	// Examples include "stop" (end of generation) or "length" (max tokens reached).
	finish_reason string

	// index is the position of this choice in the list of completions.
	index int

	// message is the generated message for this choice.
	// It contains the content and role of the response.
	message ChatCompletionMessage
}

// Usage provides details about token usage for a chat completion request.
// It includes counts for prompt, completion, and total tokens.
pub struct Usage {
pub:
	// completion_tokens is the number of tokens used in the generated response.
	completion_tokens int

	// prompt_tokens is the number of tokens used in the input prompt.
	prompt_tokens int

	// total_tokens is the total number of tokens used in the request and response.
	// This is the sum of completion_tokens and prompt_tokens.
	total_tokens int
}

// ChatCompletionResponse represents the response from the chat completion API.
// It includes the generated choices, metadata, and token usage information.
pub struct ChatCompletionResponse {
pub:
	// choices is a list of choices generated by the model.
	// Each choice includes a generated message and its associated metadata.
	choices []Choice

	// created is a Unix timestamp indicating when the response was created.
	created i64

	// id is a unique identifier for the response.
	id string

	// model specifies the name of the model used for the chat completion.
	model string

	// object is the type of object represented by this response.
	// Typically, this is "chat.completion".
	object string

	// system_fingerprint is a unique fingerprint for the system handling the request.
	system_fingerprint string

	// usage provides details about the token usage for the request and response.
	usage Usage
}

// new creates a new instance of ChatCompletionInput.
//
// Parameters:
// - messages: A list of ChatCompletionMessage objects representing the conversation history.
// - model: The name of the model to use for generating the chat completion.
//
// Returns:
// - A new instance of ChatCompletionInput.
//
// Example:
// ```v
// messages := [
//     ChatCompletionMessage{
//         role: 'user'
//         content: 'Hello!'
//     }
// ]
// input := ChatCompletionInput.new(messages, 'grok-beta')
// println(input)
// ```
pub fn ChatCompletionInput.new(messages []ChatCompletionMessage, model string) ChatCompletionInput {
	return ChatCompletionInput{
		messages: messages
		model:    model
	}
}

// get_chat_completion sends a chat completion request to the X.AI API and retrieves the response.
//
// Parameters:
// - input: A ChatCompletionInput struct containing the messages and model information for the request.
//
// Returns:
// - A ChatCompletionResponse struct containing the generated chat completion and metadata.
// - An error if the request fails or the response cannot be decoded.
//
// Example:
// ```v
// messages := [
//     ChatCompletionMessage{
//         role: 'user'
//         content: 'Tell me a joke!'
//     }
// ]
// input := ChatCompletionInput.new(messages, 'grok-beta')
// response := client.get_chat_completion(input) or { panic(err) }
// println('Generated Response: ${response.choices[0].message.content}')
// ```
pub fn (c XAIClient) get_chat_completion(input ChatCompletionInput) !ChatCompletionResponse {
	data := json.encode(input)
	res := c.post('chat/completions', data) or { return error('Failed to post chat completion') }
	return json.decode(ChatCompletionResponse, res.body) or {
		return error('Failed to decode response')
	}
}
