module vxai

import json

// The API path for language models.
pub const language_model_path = 'language-models'

// LanguageModel represents a specific language model available in the X.AI API.
// It includes details about the model's ID, creation time, input/output capabilities, and pricing.
pub struct LanguageModel {
pub:
	// completion_text_token_price specifies the token price for text completions generated by the model.
	completion_text_token_price i64

	// created is the Unix timestamp indicating when the model was created.
	created i64

	// id is the unique identifier for the language model.
	id string

	// input_modalities lists the types of input supported by the model, such as "text" or "image".
	input_modalities []string

	// object specifies the type of object represented, typically "model".
	object string

	// output_modalities lists the types of output that the model can generate, such as "text".
	output_modalities []string

	// owned_by indicates the owner of the model, usually the organization or team responsible for it.
	owned_by string

	// prompt_image_token_price specifies the token price for image-based inputs.
	prompt_image_token_price i64

	// prompt_text_token_price specifies the token price for text-based inputs.
	prompt_text_token_price i64
}

// LanguageModelsResponse represents the response from the API when querying for all available language models.
// It contains a list of LanguageModel objects.
pub struct LanguageModelsResponse {
pub:
	// models is the list of language models available in the API.
	models []LanguageModel
}

// get_language_models retrieves all available language models from the X.AI API.
//
// Returns:
// - A LanguageModelsResponse struct containing a list of all available language models.
// - An error if the request fails or if the response cannot be decoded.
pub fn (c XAIClient) get_language_models() !LanguageModelsResponse {
	res := c.get(vxai.language_model_path) or { return error('Failed to get language models') }
	return json.decode(LanguageModelsResponse, res.body) or {
		return error('Failed to decode response')
	}
}

// get_language_model retrieves details about a specific language model by its ID.
//
// Parameters:
// - id: The unique identifier of the language model to retrieve.
//
// Returns:
// - A LanguageModel struct containing details about the requested model.
// - An error if the request fails or if the response cannot be decoded.
pub fn (c XAIClient) get_language_model(id string) !LanguageModel {
	res := c.get(vxai.language_model_path + '/' + id) or { return error('Failed to get language model') }
	return json.decode(LanguageModel, res.body) or { return error('Failed to decode response') }
}
